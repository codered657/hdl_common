--  Trigonometry Package
--
--  Description: This package contains trigonometric functions and constants.
--
--  Notes: None.
--
--  Revision History:
--      Steven Okai     07/26/14    1) Initial revision.
--

library ieee;
use ieee.std_logic_1164.all;
use work.GeneralFuncPkg.all;

package TrigPkg is
    constant SINE_2048  : slv_32_vector(0 to 1023);

end TrigPkg;

package body TrigPkg is
    constant SINE_2048  : slv_32_vector(0 to 1023) := (
        x"00000000", x"006487e2", x"00c90f87", x"012d96b0", x"01921d1f", x"01f6a296", x"025b26d7", x"02bfa9a4", 
        x"03242abe", x"0388a9e9", x"03ed26e6", x"0451a176", x"04b6195d", x"051a8e5b", x"057f0034", x"05e36ea9", 
        x"0647d97c", x"06ac406f", x"0710a344", x"077501be", x"07d95b9e", x"083db0a7", x"08a2009a", x"09064b3a", 
        x"096a9049", x"09cecf89", x"0a3308bc", x"0a973ba5", x"0afb6805", x"0b5f8d9f", x"0bc3ac35", x"0c27c389", 
        x"0c8bd35e", x"0cefdb75", x"0d53db92", x"0db7d376", x"0e1bc2e3", x"0e7fa99d", x"0ee38765", x"0f475bfe", 
        x"0fab272b", x"100ee8ad", x"1072a047", x"10d64dbc", x"1139f0ce", x"119d8940", x"120116d4", x"1264994d", 
        x"12c8106e", x"132b7bf9", x"138edbb0", x"13f22f57", x"145576b1", x"14b8b17f", x"151bdf85", x"157f0086", 
        x"15e21444", x"16451a83", x"16a81304", x"170afd8d", x"176dd9de", x"17d0a7bb", x"183366e8", x"18961727", 
        x"18f8b83c", x"195b49e9", x"19bdcbf2", x"1a203e1b", x"1a82a025", x"1ae4f1d5", x"1b4732ef", x"1ba96334", 
        x"1c0b826a", x"1c6d9053", x"1ccf8cb3", x"1d31774d", x"1d934fe5", x"1df5163f", x"1e56ca1e", x"1eb86b46", 
        x"1f19f97b", x"1f7b7480", x"1fdcdc1a", x"203e300d", x"209f701c", x"21009c0b", x"2161b39f", x"21c2b69c", 
        x"2223a4c5", x"22847ddf", x"22e541ae", x"2345eff7", x"23a6887e", x"24070b07", x"24677757", x"24c7cd32", 
        x"25280c5d", x"2588349d", x"25e845b5", x"26483f6c", x"26a82185", x"2707ebc6", x"27679df4", x"27c737d2", 
        x"2826b928", x"288621b9", x"28e5714a", x"2944a7a2", x"29a3c484", x"2a02c7b8", x"2a61b101", x"2ac08025", 
        x"2b1f34eb", x"2b7dcf17", x"2bdc4e6f", x"2c3ab2b9", x"2c98fbba", x"2cf72939", x"2d553afb", x"2db330c7", 
        x"2e110a61", x"2e6ec792", x"2ecc681e", x"2f29ebcc", x"2f875262", x"2fe49ba6", x"3041c760", x"309ed555", 
        x"30fbc54d", x"3158970d", x"31b54a5d", x"3211df03", x"326e54c7", x"32caab6f", x"3326e2c2", x"3382fa88", 
        x"33def287", x"343aca87", x"3496824f", x"34f219a7", x"354d9056", x"35a8e624", x"36041ad8", x"365f2e3b", 
        x"36ba2013", x"3714f029", x"376f9e46", x"37ca2a2f", x"382493b0", x"387eda8e", x"38d8fe93", x"3932ff87", 
        x"398cdd32", x"39e6975d", x"3a402dd1", x"3a99a057", x"3af2eeb7", x"3b4c18b9", x"3ba51e29", x"3bfdfecd", 
        x"3c56ba70", x"3caf50da", x"3d07c1d5", x"3d600d2b", x"3db832a5", x"3e10320d", x"3e680b2c", x"3ebfbdcc", 
        x"3f1749b7", x"3f6eaeb8", x"3fc5ec97", x"401d0320", x"4073f21d", x"40cab957", x"4121589a", x"4177cfb0", 
        x"41ce1e64", x"42244480", x"427a41d0", x"42d0161e", x"4325c135", x"437b42e1", x"43d09aec", x"4425c923", 
        x"447acd50", x"44cfa73f", x"452456bc", x"4578db93", x"45cd358f", x"4621647c", x"46756827", x"46c9405c", 
        x"471cece6", x"47706d93", x"47c3c22e", x"4816ea85", x"4869e664", x"48bcb598", x"490f57ee", x"4961cd32", 
        x"49b41533", x"4a062fbd", x"4a581c9d", x"4aa9dba1", x"4afb6c97", x"4b4ccf4d", x"4b9e038f", x"4bef092d", 
        x"4c3fdff3", x"4c9087b1", x"4ce10034", x"4d31494b", x"4d8162c4", x"4dd14c6e", x"4e210617", x"4e708f8f", 
        x"4ebfe8a4", x"4f0f1126", x"4f5e08e3", x"4faccfaa", x"4ffb654d", x"5049c998", x"5097fc5e", x"50e5fd6c", 
        x"5133cc94", x"518169a4", x"51ced46e", x"521c0cc1", x"5269126e", x"52b5e545", x"53028517", x"534ef1b5", 
        x"539b2aef", x"53e73097", x"5433027d", x"547ea073", x"54ca0a4a", x"55153fd4", x"556040e2", x"55ab0d46", 
        x"55f5a4d2", x"56400757", x"568a34a9", x"56d42c99", x"571deef9", x"57677b9c", x"57b0d256", x"57f9f2f7", 
        x"5842dd54", x"588b913f", x"58d40e8c", x"591c550d", x"59646497", x"59ac3cfd", x"59f3de12", x"5a3b47aa", 
        x"5a827999", x"5ac973b4", x"5b1035cf", x"5b56bfbd", x"5b9d1153", x"5be32a67", x"5c290acc", x"5c6eb258", 
        x"5cb420df", x"5cf95638", x"5d3e5236", x"5d8314b0", x"5dc79d7c", x"5e0bec6e", x"5e50015d", x"5e93dc1e", 
        x"5ed77c89", x"5f1ae273", x"5f5e0db3", x"5fa0fe1e", x"5fe3b38d", x"60262dd5", x"60686cce", x"60aa704f", 
        x"60ec382f", x"612dc446", x"616f146b", x"61b02876", x"61f1003e", x"62319b9d", x"6271fa69", x"62b21c7b", 
        x"62f201ac", x"6331a9d4", x"637114cc", x"63b0426d", x"63ef328f", x"642de50d", x"646c59bf", x"64aa907f", 
        x"64e88926", x"6526438e", x"6563bf92", x"65a0fd0a", x"65ddfbd3", x"661abbc5", x"66573cbb", x"66937e90", 
        x"66cf811f", x"670b4443", x"6746c7d7", x"67820bb6", x"67bd0fbc", x"67f7d3c4", x"683257aa", x"686c9b4b", 
        x"68a69e81", x"68e06129", x"6919e320", x"69532442", x"698c246c", x"69c4e37a", x"69fd614a", x"6a359db9", 
        x"6a6d98a4", x"6aa551e8", x"6adcc964", x"6b13fef4", x"6b4af278", x"6b81a3cd", x"6bb812d0", x"6bee3f62", 
        x"6c242960", x"6c59d0a9", x"6c8f351c", x"6cc45697", x"6cf934fb", x"6d2dd027", x"6d6227fa", x"6d963c53", 
        x"6dca0d14", x"6dfd9a1b", x"6e30e349", x"6e63e87f", x"6e96a99c", x"6ec92682", x"6efb5f12", x"6f2d532c", 
        x"6f5f02b1", x"6f906d84", x"6fc19385", x"6ff27496", x"70231099", x"70536771", x"708378fe", x"70b34524", 
        x"70e2cbc6", x"71120cc5", x"71410804", x"716fbd67", x"719e2cd2", x"71cc5626", x"71fa3948", x"7227d61c", 
        x"72552c84", x"72823c66", x"72af05a6", x"72db8828", x"7307c3cf", x"7333b883", x"735f6626", x"738acc9e", 
        x"73b5ebd0", x"73e0c3a3", x"740b53fa", x"74359cbd", x"745f9dd0", x"7489571b", x"74b2c883", x"74dbf1ef", 
        x"7504d345", x"752d6c6c", x"7555bd4b", x"757dc5ca", x"75a585cf", x"75ccfd42", x"75f42c0a", x"761b1211", 
        x"7641af3c", x"76680376", x"768e0ea5", x"76b3d0b3", x"76d94988", x"76fe790e", x"77235f2d", x"7747fbce", 
        x"776c4edb", x"7790583d", x"77b417df", x"77d78daa", x"77fab988", x"781d9b64", x"78403328", x"786280bf", 
        x"78848413", x"78a63d10", x"78c7aba1", x"78e8cfb1", x"7909a92c", x"792a37fe", x"794a7c11", x"796a7554", 
        x"798a23b1", x"79a98715", x"79c89f6d", x"79e76ca6", x"7a05eead", x"7a24256e", x"7a4210d8", x"7a5fb0d8", 
        x"7a7d055b", x"7a9a0e4f", x"7ab6cba3", x"7ad33d45", x"7aef6323", x"7b0b3d2c", x"7b26cb4f", x"7b420d7a", 
        x"7b5d039d", x"7b77ada8", x"7b920b89", x"7bac1d31", x"7bc5e28f", x"7bdf5b94", x"7bf88830", x"7c116853", 
        x"7c29fbee", x"7c4242f2", x"7c5a3d4f", x"7c71eaf8", x"7c894bdd", x"7ca05ff1", x"7cb72724", x"7ccda168", 
        x"7ce3ceb1", x"7cf9aef0", x"7d0f4217", x"7d24881a", x"7d3980ec", x"7d4e2c7e", x"7d628ac5", x"7d769bb5", 
        x"7d8a5f3f", x"7d9dd55a", x"7db0fdf7", x"7dc3d90d", x"7dd6668e", x"7de8a670", x"7dfa98a7", x"7e0c3d29", 
        x"7e1d93e9", x"7e2e9cdf", x"7e3f57fe", x"7e4fc53e", x"7e5fe493", x"7e6fb5f3", x"7e7f3956", x"7e8e6eb1", 
        x"7e9d55fc", x"7eabef2c", x"7eba3a39", x"7ec8371a", x"7ed5e5c6", x"7ee34635", x"7ef0585f", x"7efd1c3c", 
        x"7f0991c3", x"7f15b8ed", x"7f2191b3", x"7f2d1c0e", x"7f3857f5", x"7f434563", x"7f4de450", x"7f5834b6", 
        x"7f62368f", x"7f6be9d4", x"7f754e7f", x"7f7e648b", x"7f872bf2", x"7f8fa4af", x"7f97cebc", x"7f9faa15", 
        x"7fa736b4", x"7fae7494", x"7fb563b2", x"7fbc040a", x"7fc25596", x"7fc85853", x"7fce0c3e", x"7fd37152", 
        x"7fd8878d", x"7fdd4eec", x"7fe1c76b", x"7fe5f108", x"7fe9cbbf", x"7fed5790", x"7ff09477", x"7ff38273", 
        x"7ff62182", x"7ff871a1", x"7ffa72d1", x"7ffc250f", x"7ffd885a", x"7ffe9cb2", x"7fff6216", x"7fffd885", 
        x"7fffffff", x"7fffd885", x"7fff6216", x"7ffe9cb2", x"7ffd885a", x"7ffc250f", x"7ffa72d1", x"7ff871a1", 
        x"7ff62182", x"7ff38273", x"7ff09477", x"7fed5790", x"7fe9cbbf", x"7fe5f108", x"7fe1c76b", x"7fdd4eec", 
        x"7fd8878d", x"7fd37152", x"7fce0c3e", x"7fc85853", x"7fc25596", x"7fbc040a", x"7fb563b2", x"7fae7494", 
        x"7fa736b4", x"7f9faa15", x"7f97cebc", x"7f8fa4af", x"7f872bf2", x"7f7e648b", x"7f754e7f", x"7f6be9d4", 
        x"7f62368f", x"7f5834b6", x"7f4de450", x"7f434563", x"7f3857f5", x"7f2d1c0e", x"7f2191b3", x"7f15b8ed", 
        x"7f0991c3", x"7efd1c3c", x"7ef0585f", x"7ee34635", x"7ed5e5c6", x"7ec8371a", x"7eba3a39", x"7eabef2c", 
        x"7e9d55fc", x"7e8e6eb1", x"7e7f3956", x"7e6fb5f3", x"7e5fe493", x"7e4fc53e", x"7e3f57fe", x"7e2e9cdf", 
        x"7e1d93e9", x"7e0c3d29", x"7dfa98a7", x"7de8a670", x"7dd6668e", x"7dc3d90d", x"7db0fdf7", x"7d9dd55a", 
        x"7d8a5f3f", x"7d769bb5", x"7d628ac5", x"7d4e2c7e", x"7d3980ec", x"7d24881a", x"7d0f4217", x"7cf9aef0", 
        x"7ce3ceb1", x"7ccda168", x"7cb72724", x"7ca05ff1", x"7c894bdd", x"7c71eaf8", x"7c5a3d4f", x"7c4242f2", 
        x"7c29fbee", x"7c116853", x"7bf88830", x"7bdf5b94", x"7bc5e28f", x"7bac1d31", x"7b920b89", x"7b77ada8", 
        x"7b5d039d", x"7b420d7a", x"7b26cb4f", x"7b0b3d2c", x"7aef6323", x"7ad33d45", x"7ab6cba3", x"7a9a0e4f", 
        x"7a7d055b", x"7a5fb0d8", x"7a4210d8", x"7a24256e", x"7a05eead", x"79e76ca6", x"79c89f6d", x"79a98715", 
        x"798a23b1", x"796a7554", x"794a7c11", x"792a37fe", x"7909a92c", x"78e8cfb1", x"78c7aba1", x"78a63d10", 
        x"78848413", x"786280bf", x"78403328", x"781d9b64", x"77fab988", x"77d78daa", x"77b417df", x"7790583d", 
        x"776c4edb", x"7747fbce", x"77235f2d", x"76fe790e", x"76d94988", x"76b3d0b3", x"768e0ea5", x"76680376", 
        x"7641af3c", x"761b1211", x"75f42c0a", x"75ccfd42", x"75a585cf", x"757dc5ca", x"7555bd4b", x"752d6c6c", 
        x"7504d345", x"74dbf1ef", x"74b2c883", x"7489571b", x"745f9dd0", x"74359cbd", x"740b53fa", x"73e0c3a3", 
        x"73b5ebd0", x"738acc9e", x"735f6626", x"7333b883", x"7307c3cf", x"72db8828", x"72af05a6", x"72823c66", 
        x"72552c84", x"7227d61c", x"71fa3948", x"71cc5626", x"719e2cd2", x"716fbd67", x"71410804", x"71120cc5", 
        x"70e2cbc6", x"70b34524", x"708378fe", x"70536771", x"70231099", x"6ff27496", x"6fc19385", x"6f906d84", 
        x"6f5f02b1", x"6f2d532c", x"6efb5f12", x"6ec92682", x"6e96a99c", x"6e63e87f", x"6e30e349", x"6dfd9a1b", 
        x"6dca0d14", x"6d963c53", x"6d6227fa", x"6d2dd027", x"6cf934fb", x"6cc45697", x"6c8f351c", x"6c59d0a9", 
        x"6c242960", x"6bee3f62", x"6bb812d0", x"6b81a3cd", x"6b4af278", x"6b13fef4", x"6adcc964", x"6aa551e8", 
        x"6a6d98a4", x"6a359db9", x"69fd614a", x"69c4e37a", x"698c246c", x"69532442", x"6919e320", x"68e06129", 
        x"68a69e81", x"686c9b4b", x"683257aa", x"67f7d3c4", x"67bd0fbc", x"67820bb6", x"6746c7d7", x"670b4443", 
        x"66cf811f", x"66937e90", x"66573cbb", x"661abbc5", x"65ddfbd3", x"65a0fd0a", x"6563bf92", x"6526438e", 
        x"64e88926", x"64aa907f", x"646c59bf", x"642de50d", x"63ef328f", x"63b0426d", x"637114cc", x"6331a9d4", 
        x"62f201ac", x"62b21c7b", x"6271fa69", x"62319b9d", x"61f1003e", x"61b02876", x"616f146b", x"612dc446", 
        x"60ec382f", x"60aa704f", x"60686cce", x"60262dd5", x"5fe3b38d", x"5fa0fe1e", x"5f5e0db3", x"5f1ae273", 
        x"5ed77c89", x"5e93dc1e", x"5e50015d", x"5e0bec6e", x"5dc79d7c", x"5d8314b0", x"5d3e5236", x"5cf95638", 
        x"5cb420df", x"5c6eb258", x"5c290acc", x"5be32a67", x"5b9d1153", x"5b56bfbd", x"5b1035cf", x"5ac973b4", 
        x"5a827999", x"5a3b47aa", x"59f3de12", x"59ac3cfd", x"59646497", x"591c550d", x"58d40e8c", x"588b913f", 
        x"5842dd54", x"57f9f2f7", x"57b0d256", x"57677b9c", x"571deef9", x"56d42c99", x"568a34a9", x"56400757", 
        x"55f5a4d2", x"55ab0d46", x"556040e2", x"55153fd4", x"54ca0a4a", x"547ea073", x"5433027d", x"53e73097", 
        x"539b2aef", x"534ef1b5", x"53028517", x"52b5e545", x"5269126e", x"521c0cc1", x"51ced46e", x"518169a4", 
        x"5133cc94", x"50e5fd6c", x"5097fc5e", x"5049c998", x"4ffb654d", x"4faccfaa", x"4f5e08e3", x"4f0f1126", 
        x"4ebfe8a4", x"4e708f8f", x"4e210617", x"4dd14c6e", x"4d8162c4", x"4d31494b", x"4ce10034", x"4c9087b1", 
        x"4c3fdff3", x"4bef092d", x"4b9e038f", x"4b4ccf4d", x"4afb6c97", x"4aa9dba1", x"4a581c9d", x"4a062fbd", 
        x"49b41533", x"4961cd32", x"490f57ee", x"48bcb598", x"4869e664", x"4816ea85", x"47c3c22e", x"47706d93", 
        x"471cece6", x"46c9405c", x"46756827", x"4621647c", x"45cd358f", x"4578db93", x"452456bc", x"44cfa73f", 
        x"447acd50", x"4425c923", x"43d09aec", x"437b42e1", x"4325c135", x"42d0161e", x"427a41d0", x"42244480", 
        x"41ce1e64", x"4177cfb0", x"4121589a", x"40cab957", x"4073f21d", x"401d0320", x"3fc5ec97", x"3f6eaeb8", 
        x"3f1749b7", x"3ebfbdcc", x"3e680b2c", x"3e10320d", x"3db832a5", x"3d600d2b", x"3d07c1d5", x"3caf50da", 
        x"3c56ba70", x"3bfdfecd", x"3ba51e29", x"3b4c18b9", x"3af2eeb7", x"3a99a057", x"3a402dd1", x"39e6975d", 
        x"398cdd32", x"3932ff87", x"38d8fe93", x"387eda8e", x"382493b0", x"37ca2a2f", x"376f9e46", x"3714f029", 
        x"36ba2013", x"365f2e3b", x"36041ad8", x"35a8e624", x"354d9056", x"34f219a7", x"3496824f", x"343aca87", 
        x"33def287", x"3382fa88", x"3326e2c2", x"32caab6f", x"326e54c7", x"3211df03", x"31b54a5d", x"3158970d", 
        x"30fbc54d", x"309ed555", x"3041c760", x"2fe49ba6", x"2f875262", x"2f29ebcc", x"2ecc681e", x"2e6ec792", 
        x"2e110a61", x"2db330c7", x"2d553afb", x"2cf72939", x"2c98fbba", x"2c3ab2b9", x"2bdc4e6f", x"2b7dcf17", 
        x"2b1f34eb", x"2ac08025", x"2a61b101", x"2a02c7b8", x"29a3c484", x"2944a7a2", x"28e5714a", x"288621b9", 
        x"2826b928", x"27c737d2", x"27679df4", x"2707ebc6", x"26a82185", x"26483f6c", x"25e845b5", x"2588349d", 
        x"25280c5d", x"24c7cd32", x"24677757", x"24070b07", x"23a6887e", x"2345eff7", x"22e541ae", x"22847ddf", 
        x"2223a4c5", x"21c2b69c", x"2161b39f", x"21009c0b", x"209f701c", x"203e300d", x"1fdcdc1a", x"1f7b7480", 
        x"1f19f97b", x"1eb86b46", x"1e56ca1e", x"1df5163f", x"1d934fe5", x"1d31774d", x"1ccf8cb3", x"1c6d9053", 
        x"1c0b826a", x"1ba96334", x"1b4732ef", x"1ae4f1d5", x"1a82a025", x"1a203e1b", x"19bdcbf2", x"195b49e9", 
        x"18f8b83c", x"18961727", x"183366e8", x"17d0a7bb", x"176dd9de", x"170afd8d", x"16a81304", x"16451a83", 
        x"15e21444", x"157f0086", x"151bdf85", x"14b8b17f", x"145576b1", x"13f22f57", x"138edbb0", x"132b7bf9", 
        x"12c8106e", x"1264994d", x"120116d4", x"119d8940", x"1139f0ce", x"10d64dbc", x"1072a047", x"100ee8ad", 
        x"0fab272b", x"0f475bfe", x"0ee38765", x"0e7fa99d", x"0e1bc2e3", x"0db7d376", x"0d53db92", x"0cefdb75", 
        x"0c8bd35e", x"0c27c389", x"0bc3ac35", x"0b5f8d9f", x"0afb6805", x"0a973ba5", x"0a3308bc", x"09cecf89", 
        x"096a9049", x"09064b3a", x"08a2009a", x"083db0a7", x"07d95b9e", x"077501be", x"0710a344", x"06ac406f", 
        x"0647d97c", x"05e36ea9", x"057f0034", x"051a8e5b", x"04b6195d", x"0451a176", x"03ed26e6", x"0388a9e9", 
        x"03242abe", x"02bfa9a4", x"025b26d7", x"01f6a296", x"01921d1f", x"012d96b0", x"00c90f87", x"006487e2");
        
end TrigPkg;